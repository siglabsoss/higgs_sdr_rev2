// don't include this file for higgs3 for now
`define LMK04133_CFG_PATH "../ti_cfg_rom_files/lmk04133_cfg_rom_ti_code_loader_950.hex"